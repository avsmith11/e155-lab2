// Avery Smith, 9/8/24, avsmith@hmc.edu
// adds 2 4-bit numbers and outputs an active low 5-bit sum
module adder(input logic [3:0] s1, s2,
			  output logic [4:0] sum
);
	assign sum = s1+s2;
endmodule
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
// putting this here so this file is for more than one line of verilog :|
